//==================================================
// Author : Tejas-Academy
// Email  : info@tejas-academy.com
// Date   : 22-03-2025
//==================================================
`include "uart_ip_tb.sv"
`include "uart_base_test.sv"
`include "uart_rdwr_test.sv"
